module seven_seg_scanner(
    input div_clock,
    input reset,
    output [3:0] anode
);

endmodule